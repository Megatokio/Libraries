/*
	this file is included by index.cgi
*/


var TITLE = «Variables class Var»
var DESCRIPTION = «c++ class for Variables in interpreter languages.»
var KEYWORDS =    «vipsi, vip script, variables, c++»
var ROBOTS = «index,nofollow»



var MAIN = 
«
h4	c++ class Var.
p	This class implements variables for interpreter languages. Basic types are number, text, list and procedure.
p	This version is currently under heavy rework. Please get the <a href="../var.stable">stable version</a> instead.
»
